/*****************************************
    
    Team XX : 
        2024000000    Kim Mina
        2024000001    Lee Minho
*****************************************/



////////////////////////////////////
//  TOP MODULE
////////////////////////////////////
module macarray (
	input CLK, RSTN, START,
	input	[11:0] MNT,
	
	output EN_I,
	output[3:0] ADDR_I,
	input [31:0] RDATA_I,
	
	output EN_W,
	output [3:0] ADDR_W,
	input [31:0] RDATA_W,

	output EN_O, RW_O,
	output [3:0] ADDR_O,
	output [63:0] WDATA_O,
	input [63:0] RDATA_O
);


	// WRITE YOUR CONTROL SYSTEM CODE




	// WRITE YOUR MAC_ARRAY DATAPATH CODE
	


endmodule
